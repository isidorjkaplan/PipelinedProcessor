module dct_rom(output logic signed [15:0] cos_q15[64]);
	assign cos_q15[0] = 32767;
	assign cos_q15[1] = 32610;
	assign cos_q15[2] = 32138;
	assign cos_q15[3] = 31357;
	assign cos_q15[4] = 30273;
	assign cos_q15[5] = 28898;
	assign cos_q15[6] = 27245;
	assign cos_q15[7] = 25330;
	assign cos_q15[8] = 23170;
	assign cos_q15[9] = 20787;
	assign cos_q15[10] = 18204;
	assign cos_q15[11] = 15446;
	assign cos_q15[12] = 12539;
	assign cos_q15[13] = 9512;
	assign cos_q15[14] = 6392;
	assign cos_q15[15] = 3211;
	assign cos_q15[16] = 0;
	assign cos_q15[17] = -3211;
	assign cos_q15[18] = -6392;
	assign cos_q15[19] = -9512;
	assign cos_q15[20] = -12539;
	assign cos_q15[21] = -15446;
	assign cos_q15[22] = -18204;
	assign cos_q15[23] = -20787;
	assign cos_q15[24] = -23170;
	assign cos_q15[25] = -25330;
	assign cos_q15[26] = -27245;
	assign cos_q15[27] = -28898;
	assign cos_q15[28] = -30273;
	assign cos_q15[29] = -31357;
	assign cos_q15[30] = -32138;
	assign cos_q15[31] = -32610;
	assign cos_q15[32] = -32768;
	assign cos_q15[33] = -32610;
	assign cos_q15[34] = -32138;
	assign cos_q15[35] = -31357;
	assign cos_q15[36] = -30273;
	assign cos_q15[37] = -28898;
	assign cos_q15[38] = -27245;
	assign cos_q15[39] = -25330;
	assign cos_q15[40] = -23170;
	assign cos_q15[41] = -20787;
	assign cos_q15[42] = -18204;
	assign cos_q15[43] = -15446;
	assign cos_q15[44] = -12539;
	assign cos_q15[45] = -9512;
	assign cos_q15[46] = -6392;
	assign cos_q15[47] = -3211;
	assign cos_q15[48] = 0;
	assign cos_q15[49] = 3211;
	assign cos_q15[50] = 6392;
	assign cos_q15[51] = 9512;
	assign cos_q15[52] = 12539;
	assign cos_q15[53] = 15446;
	assign cos_q15[54] = 18204;
	assign cos_q15[55] = 20787;
	assign cos_q15[56] = 23170;
	assign cos_q15[57] = 25330;
	assign cos_q15[58] = 27245;
	assign cos_q15[59] = 28898;
	assign cos_q15[60] = 30273;
	assign cos_q15[61] = 31357;
	assign cos_q15[62] = 32138;
	assign cos_q15[63] = 32610;
endmodule
