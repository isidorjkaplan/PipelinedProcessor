module dct_rom(output logic signed [15:0] cos_q15[129]);
	assign cos_q15[0] = 32767;
	assign cos_q15[1] = 32758;
	assign cos_q15[2] = 32728;
	assign cos_q15[3] = 32679;
	assign cos_q15[4] = 32610;
	assign cos_q15[5] = 32521;
	assign cos_q15[6] = 32413;
	assign cos_q15[7] = 32285;
	assign cos_q15[8] = 32138;
	assign cos_q15[9] = 31971;
	assign cos_q15[10] = 31785;
	assign cos_q15[11] = 31581;
	assign cos_q15[12] = 31357;
	assign cos_q15[13] = 31114;
	assign cos_q15[14] = 30852;
	assign cos_q15[15] = 30572;
	assign cos_q15[16] = 30273;
	assign cos_q15[17] = 29956;
	assign cos_q15[18] = 29621;
	assign cos_q15[19] = 29269;
	assign cos_q15[20] = 28898;
	assign cos_q15[21] = 28511;
	assign cos_q15[22] = 28106;
	assign cos_q15[23] = 27684;
	assign cos_q15[24] = 27245;
	assign cos_q15[25] = 26790;
	assign cos_q15[26] = 26319;
	assign cos_q15[27] = 25832;
	assign cos_q15[28] = 25330;
	assign cos_q15[29] = 24812;
	assign cos_q15[30] = 24279;
	assign cos_q15[31] = 23732;
	assign cos_q15[32] = 23170;
	assign cos_q15[33] = 22594;
	assign cos_q15[34] = 22005;
	assign cos_q15[35] = 21403;
	assign cos_q15[36] = 20787;
	assign cos_q15[37] = 20159;
	assign cos_q15[38] = 19519;
	assign cos_q15[39] = 18868;
	assign cos_q15[40] = 18204;
	assign cos_q15[41] = 17530;
	assign cos_q15[42] = 16846;
	assign cos_q15[43] = 16151;
	assign cos_q15[44] = 15446;
	assign cos_q15[45] = 14732;
	assign cos_q15[46] = 14010;
	assign cos_q15[47] = 13278;
	assign cos_q15[48] = 12539;
	assign cos_q15[49] = 11793;
	assign cos_q15[50] = 11039;
	assign cos_q15[51] = 10278;
	assign cos_q15[52] = 9512;
	assign cos_q15[53] = 8739;
	assign cos_q15[54] = 7961;
	assign cos_q15[55] = 7179;
	assign cos_q15[56] = 6392;
	assign cos_q15[57] = 5602;
	assign cos_q15[58] = 4808;
	assign cos_q15[59] = 4011;
	assign cos_q15[60] = 3211;
	assign cos_q15[61] = 2410;
	assign cos_q15[62] = 1607;
	assign cos_q15[63] = 804;
	assign cos_q15[64] = 0;
	assign cos_q15[65] = -804;
	assign cos_q15[66] = -1607;
	assign cos_q15[67] = -2410;
	assign cos_q15[68] = -3211;
	assign cos_q15[69] = -4011;
	assign cos_q15[70] = -4808;
	assign cos_q15[71] = -5602;
	assign cos_q15[72] = -6392;
	assign cos_q15[73] = -7179;
	assign cos_q15[74] = -7961;
	assign cos_q15[75] = -8739;
	assign cos_q15[76] = -9512;
	assign cos_q15[77] = -10278;
	assign cos_q15[78] = -11039;
	assign cos_q15[79] = -11793;
	assign cos_q15[80] = -12539;
	assign cos_q15[81] = -13278;
	assign cos_q15[82] = -14010;
	assign cos_q15[83] = -14732;
	assign cos_q15[84] = -15446;
	assign cos_q15[85] = -16151;
	assign cos_q15[86] = -16846;
	assign cos_q15[87] = -17530;
	assign cos_q15[88] = -18204;
	assign cos_q15[89] = -18868;
	assign cos_q15[90] = -19519;
	assign cos_q15[91] = -20159;
	assign cos_q15[92] = -20787;
	assign cos_q15[93] = -21403;
	assign cos_q15[94] = -22005;
	assign cos_q15[95] = -22594;
	assign cos_q15[96] = -23170;
	assign cos_q15[97] = -23732;
	assign cos_q15[98] = -24279;
	assign cos_q15[99] = -24812;
	assign cos_q15[100] = -25330;
	assign cos_q15[101] = -25832;
	assign cos_q15[102] = -26319;
	assign cos_q15[103] = -26790;
	assign cos_q15[104] = -27245;
	assign cos_q15[105] = -27684;
	assign cos_q15[106] = -28106;
	assign cos_q15[107] = -28511;
	assign cos_q15[108] = -28898;
	assign cos_q15[109] = -29269;
	assign cos_q15[110] = -29621;
	assign cos_q15[111] = -29956;
	assign cos_q15[112] = -30273;
	assign cos_q15[113] = -30572;
	assign cos_q15[114] = -30852;
	assign cos_q15[115] = -31114;
	assign cos_q15[116] = -31357;
	assign cos_q15[117] = -31581;
	assign cos_q15[118] = -31785;
	assign cos_q15[119] = -31971;
	assign cos_q15[120] = -32138;
	assign cos_q15[121] = -32285;
	assign cos_q15[122] = -32413;
	assign cos_q15[123] = -32521;
	assign cos_q15[124] = -32610;
	assign cos_q15[125] = -32679;
	assign cos_q15[126] = -32728;
	assign cos_q15[127] = -32758;
	assign cos_q15[128] = -32768;
endmodule
