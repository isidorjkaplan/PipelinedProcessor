
module dct_nios (
	clk_clk);	

	input		clk_clk;
endmodule
