module dct_rom(output logic signed [15:0] cos_q15[65]);
	assign cos_q15[0] = 32767;
	assign cos_q15[1] = 32728;
	assign cos_q15[2] = 32610;
	assign cos_q15[3] = 32413;
	assign cos_q15[4] = 32138;
	assign cos_q15[5] = 31785;
	assign cos_q15[6] = 31357;
	assign cos_q15[7] = 30852;
	assign cos_q15[8] = 30273;
	assign cos_q15[9] = 29621;
	assign cos_q15[10] = 28898;
	assign cos_q15[11] = 28106;
	assign cos_q15[12] = 27245;
	assign cos_q15[13] = 26319;
	assign cos_q15[14] = 25330;
	assign cos_q15[15] = 24279;
	assign cos_q15[16] = 23170;
	assign cos_q15[17] = 22005;
	assign cos_q15[18] = 20787;
	assign cos_q15[19] = 19519;
	assign cos_q15[20] = 18204;
	assign cos_q15[21] = 16846;
	assign cos_q15[22] = 15446;
	assign cos_q15[23] = 14010;
	assign cos_q15[24] = 12539;
	assign cos_q15[25] = 11039;
	assign cos_q15[26] = 9512;
	assign cos_q15[27] = 7961;
	assign cos_q15[28] = 6392;
	assign cos_q15[29] = 4808;
	assign cos_q15[30] = 3211;
	assign cos_q15[31] = 1607;
	assign cos_q15[32] = 0;
	assign cos_q15[33] = -1607;
	assign cos_q15[34] = -3211;
	assign cos_q15[35] = -4808;
	assign cos_q15[36] = -6392;
	assign cos_q15[37] = -7961;
	assign cos_q15[38] = -9512;
	assign cos_q15[39] = -11039;
	assign cos_q15[40] = -12539;
	assign cos_q15[41] = -14010;
	assign cos_q15[42] = -15446;
	assign cos_q15[43] = -16846;
	assign cos_q15[44] = -18204;
	assign cos_q15[45] = -19519;
	assign cos_q15[46] = -20787;
	assign cos_q15[47] = -22005;
	assign cos_q15[48] = -23170;
	assign cos_q15[49] = -24279;
	assign cos_q15[50] = -25330;
	assign cos_q15[51] = -26319;
	assign cos_q15[52] = -27245;
	assign cos_q15[53] = -28106;
	assign cos_q15[54] = -28898;
	assign cos_q15[55] = -29621;
	assign cos_q15[56] = -30273;
	assign cos_q15[57] = -30852;
	assign cos_q15[58] = -31357;
	assign cos_q15[59] = -31785;
	assign cos_q15[60] = -32138;
	assign cos_q15[61] = -32413;
	assign cos_q15[62] = -32610;
	assign cos_q15[63] = -32728;
	assign cos_q15[64] = -32768;
endmodule
